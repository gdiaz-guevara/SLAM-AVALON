-- megafunction wizard: %ALTFP_DIV%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altfp_div 

-- ============================================================
-- File Name: alt_float_div.vhd
-- Megafunction Name(s):
-- 			altfp_div
--
-- Simulation Library Files(s):
-- 			
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 18.1.0 Build 625 09/12/2018 SJ Lite Edition
-- ************************************************************


--Copyright (C) 2018  Intel Corporation. All rights reserved.
--Your use of Intel Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Intel Program License 
--Subscription Agreement, the Intel Quartus Prime License Agreement,
--the Intel FPGA IP License Agreement, or other applicable license
--agreement, including, without limitation, that your use is for
--the sole purpose of programming logic devices manufactured by
--Intel and sold by Intel or its authorized distributors.  Please
--refer to the applicable agreement for further details.


--altfp_div CBX_AUTO_BLACKBOX="ALL" DENORMAL_SUPPORT="NO" DEVICE_FAMILY="Cyclone V" OPTIMIZE="AREA" PIPELINE=6 REDUCED_FUNCTIONALITY="NO" WIDTH_EXP=8 WIDTH_MAN=23 aclr clk_en clock dataa datab result
--VERSION_BEGIN 18.1 cbx_altbarrel_shift 2018:09:12:13:04:24:SJ cbx_altera_syncram_nd_impl 2018:09:12:13:04:24:SJ cbx_altfp_div 2018:09:12:13:04:24:SJ cbx_altsyncram 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_abs 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_compare 2018:09:12:13:04:24:SJ cbx_lpm_decode 2018:09:12:13:04:24:SJ cbx_lpm_divide 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_stratixiii 2018:09:12:13:04:24:SJ cbx_stratixv 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END


--altfp_div_pst CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" FILE_NAME="alt_float_div.vhd:a" PIPELINE=6 WIDTH_EXP=8 WIDTH_MAN=23 aclr clk_en clock dataa datab result
--VERSION_BEGIN 18.1 cbx_altbarrel_shift 2018:09:12:13:04:24:SJ cbx_altera_syncram_nd_impl 2018:09:12:13:04:24:SJ cbx_altfp_div 2018:09:12:13:04:24:SJ cbx_altsyncram 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_abs 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_compare 2018:09:12:13:04:24:SJ cbx_lpm_decode 2018:09:12:13:04:24:SJ cbx_lpm_divide 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_stratixiii 2018:09:12:13:04:24:SJ cbx_stratixv 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END

 LIBRARY altera_mf;
 USE altera_mf.all;

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = altsyncram 1 lpm_add_sub 4 lpm_compare 1 lpm_mult 5 mux21 74 reg 339 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  alt_float_div_altfp_div_pst_jcf IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clk_en	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC;
		 dataa	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 datab	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0)
	 ); 
 END alt_float_div_altfp_div_pst_jcf;

 ARCHITECTURE RTL OF alt_float_div_altfp_div_pst_jcf IS

	 SIGNAL  wire_altsyncram3_q_a	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL	 a_is_infinity_dffe_0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 a_is_infinity_dffe_1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_a_is_infinity_dffe_1_w_lg_q318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 a_is_infinity_dffe_2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 a_is_infinity_dffe_3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 a_is_infinity_dffe_4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 a_zero_b_not_dffe_0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 a_zero_b_not_dffe_1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_a_zero_b_not_dffe_1_w_lg_q326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 a_zero_b_not_dffe_2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 a_zero_b_not_dffe_3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 a_zero_b_not_dffe_4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 b1_dffe_0	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 b_is_infinity_dffe_0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 b_is_infinity_dffe_1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_b_is_infinity_dffe_1_w_lg_q325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 b_is_infinity_dffe_2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 b_is_infinity_dffe_3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 b_is_infinity_dffe_4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 both_exp_zeros_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 divbyzero_pipe_dffe_0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 divbyzero_pipe_dffe_1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_divbyzero_pipe_dffe_1_w_lg_q317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 divbyzero_pipe_dffe_2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 divbyzero_pipe_dffe_3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 divbyzero_pipe_dffe_4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 e1_dffe_0	:	STD_LOGIC_VECTOR(16 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 e1_dffe_1	:	STD_LOGIC_VECTOR(16 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_result_dffe_0	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_result_dffe_1	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_result_dffe_2	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_result_dffe_3	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 frac_a_smaller_dffe1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_a_dffe1_dffe1	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_b_dffe1_dffe1	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_result_dffe	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_pipe_dffe_0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_pipe_dffe_1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_nan_pipe_dffe_1_w_lg_q308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 nan_pipe_dffe_2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_pipe_dffe_3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_pipe_dffe_4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 over_under_dffe_0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 over_under_dffe_1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 over_under_dffe_2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 quotient_j_dffe	:	STD_LOGIC_VECTOR(16 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 quotient_k_dffe_0	:	STD_LOGIC_VECTOR(16 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 remainder_j_dffe_0	:	STD_LOGIC_VECTOR(49 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 remainder_j_dffe_1	:	STD_LOGIC_VECTOR(49 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_pipe_dffe_0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_pipe_dffe_1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_pipe_dffe_2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_pipe_dffe_3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_pipe_dffe_4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_pipe_dffe_5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_bias_addition_overflow	:	STD_LOGIC;
	 SIGNAL  wire_bias_addition_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_exp_sub_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_quotient_process_dataa	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_quotient_process_datab	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_quotient_process_result	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_quotient_process_w_result_range425w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_remainder_sub_0_dataa	:	STD_LOGIC_VECTOR (49 DOWNTO 0);
	 SIGNAL  wire_remainder_sub_0_result	:	STD_LOGIC_VECTOR (49 DOWNTO 0);
	 SIGNAL  wire_cmpr2_alb	:	STD_LOGIC;
	 SIGNAL  wire_a1_prod_datab	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_a1_prod_result	:	STD_LOGIC_VECTOR (34 DOWNTO 0);
	 SIGNAL  wire_b1_prod_w_lg_w_result_range358w359w	:	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  wire_b1_prod_datab	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_b1_prod_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_b1_prod_w_result_range358w	:	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  wire_q_partial_0_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_q_partial_0_w_result_range373w	:	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  wire_q_partial_1_w_lg_w_result_range407w408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_q_partial_1_w_lg_w_result_range410w411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_q_partial_1_w_lg_w_result_range413w414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_q_partial_1_w_lg_w_result_range416w417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_q_partial_1_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_q_partial_1_w_result_range407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_q_partial_1_w_result_range410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_q_partial_1_w_result_range413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_q_partial_1_w_result_range416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_remainder_mult_0_result	:	STD_LOGIC_VECTOR (50 DOWNTO 0);
	 SIGNAL	wire_exp_result_muxa_dataout	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL	wire_man_a_adjusteda_dataout	:	STD_LOGIC_VECTOR(24 DOWNTO 0);
	 SIGNAL	wire_man_result_muxa_dataout	:	STD_LOGIC_VECTOR(22 DOWNTO 0);
	 SIGNAL	wire_select_bias_2a_dataout	:	STD_LOGIC_VECTOR(8 DOWNTO 0);
	 SIGNAL	wire_select_biasa_dataout	:	STD_LOGIC_VECTOR(8 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_lg_w_lg_bias_addition_overf_w304w305w306w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_lg_bias_addition_overf_w304w305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_lg_bias_addition_overf_w304w312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w302w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_bias_addition_w_range262w285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_bias_addition_w_range265w287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_bias_addition_w_range268w289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_bias_addition_w_range271w291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_bias_addition_w_range274w293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_bias_addition_w_range277w295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_bias_addition_w_range280w297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range11w17w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range21w27w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range31w37w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range41w47w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range51w57w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range61w67w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range71w77w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range14w19w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range24w29w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range34w39w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range44w49w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range54w59w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range64w69w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range74w79w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_exp_a_all_one_w_range78w222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_exp_add_output_all_one_range298w321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_exp_b_all_one_w_range80w224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_exp_b_not_zero_w_range76w256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_a_is_infinity_w233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_a_is_nan_w234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_bias_addition_overf_w304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_exp_sign_w303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_exp_a_not_zero_w_range73w227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_man_a_not_zero_w_range215w221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_man_b_not_zero_w_range218w223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_lg_w_lg_bias_addition_overf_w299w300w301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_lg_bias_addition_overf_w299w300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_bias_addition_overf_w323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_bias_addition_overf_w299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_bias_addition_w_range262w263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_bias_addition_w_range265w266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_bias_addition_w_range268w269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_bias_addition_w_range271w272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_bias_addition_w_range274w275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_bias_addition_w_range277w278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_bias_addition_w_range280w281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range141w142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range147w148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range153w154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range159w160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range165w166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range171w172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range177w178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range183w184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range189w190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range195w196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range87w88w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range201w202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range207w208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range213w214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range11w12w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range21w22w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range31w32w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range41w42w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range51w52w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range61w62w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range93w94w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range71w72w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range99w100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range105w106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range111w112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range117w118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range123w124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range129w130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_dataa_range135w136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range144w145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range150w151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range156w157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range162w163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range168w169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range174w175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range180w181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range186w187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range192w193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range198w199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range90w91w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range204w205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range210w211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range216w217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range14w15w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range24w25w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range34w35w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range44w45w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range54w55w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range64w65w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range96w97w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range74w75w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range102w103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range108w109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range114w115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range120w121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range126w127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range132w133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_lg_w_datab_range138w139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  a_is_infinity_w :	STD_LOGIC;
	 SIGNAL  a_is_nan_w :	STD_LOGIC;
	 SIGNAL  a_zero_b_not :	STD_LOGIC;
	 SIGNAL  b1_dffe_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  b_is_infinity_w :	STD_LOGIC;
	 SIGNAL  b_is_nan_w :	STD_LOGIC;
	 SIGNAL  bias_addition_overf_w :	STD_LOGIC;
	 SIGNAL  bias_addition_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  both_exp_zeros :	STD_LOGIC;
	 SIGNAL  e0_dffe1_wo :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  e0_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  e1_w :	STD_LOGIC_VECTOR (50 DOWNTO 0);
	 SIGNAL  exp_a_all_one_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_a_not_zero_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_add_output_all_one :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_add_output_not_zero :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_b_all_one_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_b_not_zero_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_result_mux_out :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_result_mux_sel_w :	STD_LOGIC;
	 SIGNAL  exp_result_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_sign_w :	STD_LOGIC;
	 SIGNAL  exp_sub_a_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  exp_sub_b_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  exp_sub_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  frac_a_smaller_dffe1_wi :	STD_LOGIC;
	 SIGNAL  frac_a_smaller_dffe1_wo :	STD_LOGIC;
	 SIGNAL  frac_a_smaller_w :	STD_LOGIC;
	 SIGNAL  guard_bit :	STD_LOGIC;
	 SIGNAL  man_a_adjusted_w :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  man_a_dffe1_wi :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_a_dffe1_wo :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_a_not_zero_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_b_adjusted_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  man_b_dffe1_wi :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_b_dffe1_wo :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_b_not_zero_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_result_dffe_wi :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_result_dffe_wo :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_result_mux_select :	STD_LOGIC;
	 SIGNAL  man_result_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_zeros_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  overflow_ones_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  overflow_underflow :	STD_LOGIC;
	 SIGNAL  overflow_w :	STD_LOGIC;
	 SIGNAL  quotient_accumulate_w :	STD_LOGIC_VECTOR (61 DOWNTO 0);
	 SIGNAL  quotient_process_cin_w :	STD_LOGIC;
	 SIGNAL  remainder_j_w :	STD_LOGIC_VECTOR (99 DOWNTO 0);
	 SIGNAL  round_bit :	STD_LOGIC;
	 SIGNAL  select_bias_out_2_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  select_bias_out_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  sticky_bits :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  underflow_w :	STD_LOGIC;
	 SIGNAL  underflow_zeros_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  value_add_one_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  value_normal_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  value_zero_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_bias_addition_w_range262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_bias_addition_w_range265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_bias_addition_w_range268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_bias_addition_w_range271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_bias_addition_w_range274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_bias_addition_w_range277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_bias_addition_w_range280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range87w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range11w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range21w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range31w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range41w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range51w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range61w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range93w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range71w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range99w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_dataa_range135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range90w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range14w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range24w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range34w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range44w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range54w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range64w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range96w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range74w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_datab_range138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_e1_w_range360w	:	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_e1_w_range368w	:	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_a_all_one_w_range7w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_a_all_one_w_range18w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_a_all_one_w_range28w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_a_all_one_w_range38w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_a_all_one_w_range48w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_a_all_one_w_range58w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_a_all_one_w_range68w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_a_all_one_w_range78w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_a_not_zero_w_range2w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_a_not_zero_w_range13w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_a_not_zero_w_range23w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_a_not_zero_w_range33w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_a_not_zero_w_range43w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_a_not_zero_w_range53w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_a_not_zero_w_range63w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_a_not_zero_w_range73w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_add_output_all_one_range283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_add_output_all_one_range286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_add_output_all_one_range288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_add_output_all_one_range290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_add_output_all_one_range292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_add_output_all_one_range294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_add_output_all_one_range296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_add_output_all_one_range298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_add_output_not_zero_range260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_add_output_not_zero_range264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_add_output_not_zero_range267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_add_output_not_zero_range270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_add_output_not_zero_range273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_add_output_not_zero_range276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_add_output_not_zero_range279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_b_all_one_w_range9w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_b_all_one_w_range20w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_b_all_one_w_range30w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_b_all_one_w_range40w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_b_all_one_w_range50w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_b_all_one_w_range60w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_b_all_one_w_range70w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_b_all_one_w_range80w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_b_not_zero_w_range5w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_b_not_zero_w_range16w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_b_not_zero_w_range26w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_b_not_zero_w_range36w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_b_not_zero_w_range46w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_b_not_zero_w_range56w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_b_not_zero_w_range66w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_exp_b_not_zero_w_range76w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range82w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range89w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range95w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_a_not_zero_w_range137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range85w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range92w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range98w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_man_b_not_zero_w_range140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_remainder_j_w_range363w	:	STD_LOGIC_VECTOR (49 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_sticky_bits_range405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_sticky_bits_range409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_sticky_bits_range412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_sticky_bits_range415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_pst1_w_w_quotient_accumulate_w_range385w_range386w	:	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 COMPONENT  altsyncram
	 GENERIC 
	 (
		ADDRESS_ACLR_A	:	STRING := "UNUSED";
		ADDRESS_ACLR_B	:	STRING := "NONE";
		ADDRESS_REG_B	:	STRING := "CLOCK1";
		BYTE_SIZE	:	NATURAL := 8;
		BYTEENA_ACLR_A	:	STRING := "UNUSED";
		BYTEENA_ACLR_B	:	STRING := "NONE";
		BYTEENA_REG_B	:	STRING := "CLOCK1";
		CLOCK_ENABLE_CORE_A	:	STRING := "USE_INPUT_CLKEN";
		CLOCK_ENABLE_CORE_B	:	STRING := "USE_INPUT_CLKEN";
		CLOCK_ENABLE_INPUT_A	:	STRING := "NORMAL";
		CLOCK_ENABLE_INPUT_B	:	STRING := "NORMAL";
		CLOCK_ENABLE_OUTPUT_A	:	STRING := "NORMAL";
		CLOCK_ENABLE_OUTPUT_B	:	STRING := "NORMAL";
		ECC_PIPELINE_STAGE_ENABLED	:	STRING := "FALSE";
		ENABLE_ECC	:	STRING := "FALSE";
		IMPLEMENT_IN_LES	:	STRING := "OFF";
		INDATA_ACLR_A	:	STRING := "UNUSED";
		INDATA_ACLR_B	:	STRING := "NONE";
		INDATA_REG_B	:	STRING := "CLOCK1";
		INIT_FILE	:	STRING := "UNUSED";
		INIT_FILE_LAYOUT	:	STRING := "PORT_A";
		MAXIMUM_DEPTH	:	NATURAL := 0;
		NUMWORDS_A	:	NATURAL := 0;
		NUMWORDS_B	:	NATURAL := 0;
		OPERATION_MODE	:	STRING := "BIDIR_DUAL_PORT";
		OUTDATA_ACLR_A	:	STRING := "NONE";
		OUTDATA_ACLR_B	:	STRING := "NONE";
		OUTDATA_REG_A	:	STRING := "UNREGISTERED";
		OUTDATA_REG_B	:	STRING := "UNREGISTERED";
		POWER_UP_UNINITIALIZED	:	STRING := "FALSE";
		RAM_BLOCK_TYPE	:	STRING := "AUTO";
		RDCONTROL_ACLR_B	:	STRING := "NONE";
		RDCONTROL_REG_B	:	STRING := "CLOCK1";
		READ_DURING_WRITE_MODE_MIXED_PORTS	:	STRING := "DONT_CARE";
		read_during_write_mode_port_a	:	STRING := "NEW_DATA_NO_NBE_READ";
		read_during_write_mode_port_b	:	STRING := "NEW_DATA_NO_NBE_READ";
		WIDTH_A	:	NATURAL;
		WIDTH_B	:	NATURAL := 1;
		WIDTH_BYTEENA_A	:	NATURAL := 1;
		WIDTH_BYTEENA_B	:	NATURAL := 1;
		WIDTH_ECCSTATUS	:	NATURAL := 3;
		WIDTHAD_A	:	NATURAL;
		WIDTHAD_B	:	NATURAL := 1;
		WRCONTROL_ACLR_A	:	STRING := "UNUSED";
		WRCONTROL_ACLR_B	:	STRING := "NONE";
		WRCONTROL_WRADDRESS_REG_B	:	STRING := "CLOCK1";
		INTENDED_DEVICE_FAMILY	:	STRING := "Cyclone V";
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "altsyncram"
	 );
	 PORT
	 ( 
		aclr0	:	IN STD_LOGIC := '0';
		aclr1	:	IN STD_LOGIC := '0';
		address_a	:	IN STD_LOGIC_VECTOR(WIDTHAD_A-1 DOWNTO 0);
		address_b	:	IN STD_LOGIC_VECTOR(WIDTHAD_B-1 DOWNTO 0) := (OTHERS => '1');
		addressstall_a	:	IN STD_LOGIC := '0';
		addressstall_b	:	IN STD_LOGIC := '0';
		byteena_a	:	IN STD_LOGIC_VECTOR(WIDTH_BYTEENA_A-1 DOWNTO 0) := (OTHERS => '1');
		byteena_b	:	IN STD_LOGIC_VECTOR(WIDTH_BYTEENA_B-1 DOWNTO 0) := (OTHERS => '1');
		clock0	:	IN STD_LOGIC := '1';
		clock1	:	IN STD_LOGIC := '1';
		clocken0	:	IN STD_LOGIC := '1';
		clocken1	:	IN STD_LOGIC := '1';
		clocken2	:	IN STD_LOGIC := '1';
		clocken3	:	IN STD_LOGIC := '1';
		data_a	:	IN STD_LOGIC_VECTOR(WIDTH_A-1 DOWNTO 0) := (OTHERS => '1');
		data_b	:	IN STD_LOGIC_VECTOR(WIDTH_B-1 DOWNTO 0) := (OTHERS => '1');
		eccstatus	:	OUT STD_LOGIC_VECTOR(WIDTH_ECCSTATUS-1 DOWNTO 0);
		q_a	:	OUT STD_LOGIC_VECTOR(WIDTH_A-1 DOWNTO 0);
		q_b	:	OUT STD_LOGIC_VECTOR(WIDTH_B-1 DOWNTO 0);
		rden_a	:	IN STD_LOGIC := '1';
		rden_b	:	IN STD_LOGIC := '1';
		wren_a	:	IN STD_LOGIC := '0';
		wren_b	:	IN STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_mult
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTHA	:	NATURAL;
		LPM_WIDTHB	:	NATURAL;
		LPM_WIDTHP	:	NATURAL;
		LPM_WIDTHS	:	NATURAL := 1;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_mult"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTHA-1 DOWNTO 0);
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTHB-1 DOWNTO 0);
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTHP-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sum	:	IN STD_LOGIC_VECTOR(LPM_WIDTHS-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	loop0 : FOR i IN 0 TO 7 GENERATE 
		wire_altfp_div_pst1_w_lg_w_lg_w_lg_bias_addition_overf_w304w305w306w(i) <= wire_altfp_div_pst1_w_lg_w_lg_bias_addition_overf_w304w305w(0) AND bias_addition_w(i);
	END GENERATE loop0;
	wire_altfp_div_pst1_w322w(0) <= wire_altfp_div_pst1_w_lg_w_exp_add_output_all_one_range298w321w(0) AND wire_altfp_div_pst1_w_lg_exp_sign_w303w(0);
	wire_altfp_div_pst1_w_lg_w_lg_bias_addition_overf_w304w305w(0) <= wire_altfp_div_pst1_w_lg_bias_addition_overf_w304w(0) AND wire_altfp_div_pst1_w_lg_exp_sign_w303w(0);
	wire_altfp_div_pst1_w_lg_w_lg_bias_addition_overf_w304w312w(0) <= wire_altfp_div_pst1_w_lg_bias_addition_overf_w304w(0) AND exp_sign_w;
	loop1 : FOR i IN 0 TO 7 GENERATE 
		wire_altfp_div_pst1_w302w(i) <= wire_altfp_div_pst1_w_lg_w_lg_w_lg_bias_addition_overf_w299w300w301w(0) AND overflow_ones_w(i);
	END GENERATE loop1;
	wire_altfp_div_pst1_w_lg_w_bias_addition_w_range262w285w(0) <= wire_altfp_div_pst1_w_bias_addition_w_range262w(0) AND wire_altfp_div_pst1_w_exp_add_output_all_one_range283w(0);
	wire_altfp_div_pst1_w_lg_w_bias_addition_w_range265w287w(0) <= wire_altfp_div_pst1_w_bias_addition_w_range265w(0) AND wire_altfp_div_pst1_w_exp_add_output_all_one_range286w(0);
	wire_altfp_div_pst1_w_lg_w_bias_addition_w_range268w289w(0) <= wire_altfp_div_pst1_w_bias_addition_w_range268w(0) AND wire_altfp_div_pst1_w_exp_add_output_all_one_range288w(0);
	wire_altfp_div_pst1_w_lg_w_bias_addition_w_range271w291w(0) <= wire_altfp_div_pst1_w_bias_addition_w_range271w(0) AND wire_altfp_div_pst1_w_exp_add_output_all_one_range290w(0);
	wire_altfp_div_pst1_w_lg_w_bias_addition_w_range274w293w(0) <= wire_altfp_div_pst1_w_bias_addition_w_range274w(0) AND wire_altfp_div_pst1_w_exp_add_output_all_one_range292w(0);
	wire_altfp_div_pst1_w_lg_w_bias_addition_w_range277w295w(0) <= wire_altfp_div_pst1_w_bias_addition_w_range277w(0) AND wire_altfp_div_pst1_w_exp_add_output_all_one_range294w(0);
	wire_altfp_div_pst1_w_lg_w_bias_addition_w_range280w297w(0) <= wire_altfp_div_pst1_w_bias_addition_w_range280w(0) AND wire_altfp_div_pst1_w_exp_add_output_all_one_range296w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range11w17w(0) <= wire_altfp_div_pst1_w_dataa_range11w(0) AND wire_altfp_div_pst1_w_exp_a_all_one_w_range7w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range21w27w(0) <= wire_altfp_div_pst1_w_dataa_range21w(0) AND wire_altfp_div_pst1_w_exp_a_all_one_w_range18w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range31w37w(0) <= wire_altfp_div_pst1_w_dataa_range31w(0) AND wire_altfp_div_pst1_w_exp_a_all_one_w_range28w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range41w47w(0) <= wire_altfp_div_pst1_w_dataa_range41w(0) AND wire_altfp_div_pst1_w_exp_a_all_one_w_range38w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range51w57w(0) <= wire_altfp_div_pst1_w_dataa_range51w(0) AND wire_altfp_div_pst1_w_exp_a_all_one_w_range48w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range61w67w(0) <= wire_altfp_div_pst1_w_dataa_range61w(0) AND wire_altfp_div_pst1_w_exp_a_all_one_w_range58w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range71w77w(0) <= wire_altfp_div_pst1_w_dataa_range71w(0) AND wire_altfp_div_pst1_w_exp_a_all_one_w_range68w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range14w19w(0) <= wire_altfp_div_pst1_w_datab_range14w(0) AND wire_altfp_div_pst1_w_exp_b_all_one_w_range9w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range24w29w(0) <= wire_altfp_div_pst1_w_datab_range24w(0) AND wire_altfp_div_pst1_w_exp_b_all_one_w_range20w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range34w39w(0) <= wire_altfp_div_pst1_w_datab_range34w(0) AND wire_altfp_div_pst1_w_exp_b_all_one_w_range30w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range44w49w(0) <= wire_altfp_div_pst1_w_datab_range44w(0) AND wire_altfp_div_pst1_w_exp_b_all_one_w_range40w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range54w59w(0) <= wire_altfp_div_pst1_w_datab_range54w(0) AND wire_altfp_div_pst1_w_exp_b_all_one_w_range50w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range64w69w(0) <= wire_altfp_div_pst1_w_datab_range64w(0) AND wire_altfp_div_pst1_w_exp_b_all_one_w_range60w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range74w79w(0) <= wire_altfp_div_pst1_w_datab_range74w(0) AND wire_altfp_div_pst1_w_exp_b_all_one_w_range70w(0);
	wire_altfp_div_pst1_w_lg_w_exp_a_all_one_w_range78w222w(0) <= wire_altfp_div_pst1_w_exp_a_all_one_w_range78w(0) AND wire_altfp_div_pst1_w_lg_w_man_a_not_zero_w_range215w221w(0);
	wire_altfp_div_pst1_w_lg_w_exp_add_output_all_one_range298w321w(0) <= wire_altfp_div_pst1_w_exp_add_output_all_one_range298w(0) AND wire_altfp_div_pst1_w_lg_bias_addition_overf_w304w(0);
	wire_altfp_div_pst1_w_lg_w_exp_b_all_one_w_range80w224w(0) <= wire_altfp_div_pst1_w_exp_b_all_one_w_range80w(0) AND wire_altfp_div_pst1_w_lg_w_man_b_not_zero_w_range218w223w(0);
	wire_altfp_div_pst1_w_lg_w_exp_b_not_zero_w_range76w256w(0) <= wire_altfp_div_pst1_w_exp_b_not_zero_w_range76w(0) AND wire_altfp_div_pst1_w_lg_w_exp_a_not_zero_w_range73w227w(0);
	wire_altfp_div_pst1_w_lg_a_is_infinity_w233w(0) <= NOT a_is_infinity_w;
	wire_altfp_div_pst1_w_lg_a_is_nan_w234w(0) <= NOT a_is_nan_w;
	wire_altfp_div_pst1_w_lg_bias_addition_overf_w304w(0) <= NOT bias_addition_overf_w;
	wire_altfp_div_pst1_w_lg_exp_sign_w303w(0) <= NOT exp_sign_w;
	wire_altfp_div_pst1_w_lg_w_exp_a_not_zero_w_range73w227w(0) <= NOT wire_altfp_div_pst1_w_exp_a_not_zero_w_range73w(0);
	wire_altfp_div_pst1_w_lg_w_man_a_not_zero_w_range215w221w(0) <= NOT wire_altfp_div_pst1_w_man_a_not_zero_w_range215w(0);
	wire_altfp_div_pst1_w_lg_w_man_b_not_zero_w_range218w223w(0) <= NOT wire_altfp_div_pst1_w_man_b_not_zero_w_range218w(0);
	wire_altfp_div_pst1_w_lg_w_lg_w_lg_bias_addition_overf_w299w300w301w(0) <= wire_altfp_div_pst1_w_lg_w_lg_bias_addition_overf_w299w300w(0) OR a_is_infinity_dffe_1;
	wire_altfp_div_pst1_w_lg_w_lg_bias_addition_overf_w299w300w(0) <= wire_altfp_div_pst1_w_lg_bias_addition_overf_w299w(0) OR nan_pipe_dffe_1;
	wire_altfp_div_pst1_w_lg_bias_addition_overf_w323w(0) <= bias_addition_overf_w OR wire_altfp_div_pst1_w322w(0);
	wire_altfp_div_pst1_w_lg_bias_addition_overf_w299w(0) <= bias_addition_overf_w OR divbyzero_pipe_dffe_1;
	wire_altfp_div_pst1_w_lg_w_bias_addition_w_range262w263w(0) <= wire_altfp_div_pst1_w_bias_addition_w_range262w(0) OR wire_altfp_div_pst1_w_exp_add_output_not_zero_range260w(0);
	wire_altfp_div_pst1_w_lg_w_bias_addition_w_range265w266w(0) <= wire_altfp_div_pst1_w_bias_addition_w_range265w(0) OR wire_altfp_div_pst1_w_exp_add_output_not_zero_range264w(0);
	wire_altfp_div_pst1_w_lg_w_bias_addition_w_range268w269w(0) <= wire_altfp_div_pst1_w_bias_addition_w_range268w(0) OR wire_altfp_div_pst1_w_exp_add_output_not_zero_range267w(0);
	wire_altfp_div_pst1_w_lg_w_bias_addition_w_range271w272w(0) <= wire_altfp_div_pst1_w_bias_addition_w_range271w(0) OR wire_altfp_div_pst1_w_exp_add_output_not_zero_range270w(0);
	wire_altfp_div_pst1_w_lg_w_bias_addition_w_range274w275w(0) <= wire_altfp_div_pst1_w_bias_addition_w_range274w(0) OR wire_altfp_div_pst1_w_exp_add_output_not_zero_range273w(0);
	wire_altfp_div_pst1_w_lg_w_bias_addition_w_range277w278w(0) <= wire_altfp_div_pst1_w_bias_addition_w_range277w(0) OR wire_altfp_div_pst1_w_exp_add_output_not_zero_range276w(0);
	wire_altfp_div_pst1_w_lg_w_bias_addition_w_range280w281w(0) <= wire_altfp_div_pst1_w_bias_addition_w_range280w(0) OR wire_altfp_div_pst1_w_exp_add_output_not_zero_range279w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range141w142w(0) <= wire_altfp_div_pst1_w_dataa_range141w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range137w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range147w148w(0) <= wire_altfp_div_pst1_w_dataa_range147w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range143w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range153w154w(0) <= wire_altfp_div_pst1_w_dataa_range153w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range149w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range159w160w(0) <= wire_altfp_div_pst1_w_dataa_range159w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range155w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range165w166w(0) <= wire_altfp_div_pst1_w_dataa_range165w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range161w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range171w172w(0) <= wire_altfp_div_pst1_w_dataa_range171w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range167w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range177w178w(0) <= wire_altfp_div_pst1_w_dataa_range177w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range173w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range183w184w(0) <= wire_altfp_div_pst1_w_dataa_range183w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range179w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range189w190w(0) <= wire_altfp_div_pst1_w_dataa_range189w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range185w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range195w196w(0) <= wire_altfp_div_pst1_w_dataa_range195w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range191w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range87w88w(0) <= wire_altfp_div_pst1_w_dataa_range87w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range82w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range201w202w(0) <= wire_altfp_div_pst1_w_dataa_range201w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range197w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range207w208w(0) <= wire_altfp_div_pst1_w_dataa_range207w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range203w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range213w214w(0) <= wire_altfp_div_pst1_w_dataa_range213w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range209w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range11w12w(0) <= wire_altfp_div_pst1_w_dataa_range11w(0) OR wire_altfp_div_pst1_w_exp_a_not_zero_w_range2w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range21w22w(0) <= wire_altfp_div_pst1_w_dataa_range21w(0) OR wire_altfp_div_pst1_w_exp_a_not_zero_w_range13w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range31w32w(0) <= wire_altfp_div_pst1_w_dataa_range31w(0) OR wire_altfp_div_pst1_w_exp_a_not_zero_w_range23w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range41w42w(0) <= wire_altfp_div_pst1_w_dataa_range41w(0) OR wire_altfp_div_pst1_w_exp_a_not_zero_w_range33w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range51w52w(0) <= wire_altfp_div_pst1_w_dataa_range51w(0) OR wire_altfp_div_pst1_w_exp_a_not_zero_w_range43w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range61w62w(0) <= wire_altfp_div_pst1_w_dataa_range61w(0) OR wire_altfp_div_pst1_w_exp_a_not_zero_w_range53w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range93w94w(0) <= wire_altfp_div_pst1_w_dataa_range93w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range89w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range71w72w(0) <= wire_altfp_div_pst1_w_dataa_range71w(0) OR wire_altfp_div_pst1_w_exp_a_not_zero_w_range63w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range99w100w(0) <= wire_altfp_div_pst1_w_dataa_range99w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range95w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range105w106w(0) <= wire_altfp_div_pst1_w_dataa_range105w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range101w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range111w112w(0) <= wire_altfp_div_pst1_w_dataa_range111w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range107w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range117w118w(0) <= wire_altfp_div_pst1_w_dataa_range117w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range113w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range123w124w(0) <= wire_altfp_div_pst1_w_dataa_range123w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range119w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range129w130w(0) <= wire_altfp_div_pst1_w_dataa_range129w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range125w(0);
	wire_altfp_div_pst1_w_lg_w_dataa_range135w136w(0) <= wire_altfp_div_pst1_w_dataa_range135w(0) OR wire_altfp_div_pst1_w_man_a_not_zero_w_range131w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range144w145w(0) <= wire_altfp_div_pst1_w_datab_range144w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range140w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range150w151w(0) <= wire_altfp_div_pst1_w_datab_range150w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range146w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range156w157w(0) <= wire_altfp_div_pst1_w_datab_range156w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range152w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range162w163w(0) <= wire_altfp_div_pst1_w_datab_range162w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range158w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range168w169w(0) <= wire_altfp_div_pst1_w_datab_range168w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range164w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range174w175w(0) <= wire_altfp_div_pst1_w_datab_range174w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range170w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range180w181w(0) <= wire_altfp_div_pst1_w_datab_range180w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range176w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range186w187w(0) <= wire_altfp_div_pst1_w_datab_range186w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range182w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range192w193w(0) <= wire_altfp_div_pst1_w_datab_range192w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range188w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range198w199w(0) <= wire_altfp_div_pst1_w_datab_range198w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range194w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range90w91w(0) <= wire_altfp_div_pst1_w_datab_range90w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range85w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range204w205w(0) <= wire_altfp_div_pst1_w_datab_range204w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range200w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range210w211w(0) <= wire_altfp_div_pst1_w_datab_range210w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range206w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range216w217w(0) <= wire_altfp_div_pst1_w_datab_range216w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range212w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range14w15w(0) <= wire_altfp_div_pst1_w_datab_range14w(0) OR wire_altfp_div_pst1_w_exp_b_not_zero_w_range5w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range24w25w(0) <= wire_altfp_div_pst1_w_datab_range24w(0) OR wire_altfp_div_pst1_w_exp_b_not_zero_w_range16w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range34w35w(0) <= wire_altfp_div_pst1_w_datab_range34w(0) OR wire_altfp_div_pst1_w_exp_b_not_zero_w_range26w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range44w45w(0) <= wire_altfp_div_pst1_w_datab_range44w(0) OR wire_altfp_div_pst1_w_exp_b_not_zero_w_range36w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range54w55w(0) <= wire_altfp_div_pst1_w_datab_range54w(0) OR wire_altfp_div_pst1_w_exp_b_not_zero_w_range46w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range64w65w(0) <= wire_altfp_div_pst1_w_datab_range64w(0) OR wire_altfp_div_pst1_w_exp_b_not_zero_w_range56w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range96w97w(0) <= wire_altfp_div_pst1_w_datab_range96w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range92w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range74w75w(0) <= wire_altfp_div_pst1_w_datab_range74w(0) OR wire_altfp_div_pst1_w_exp_b_not_zero_w_range66w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range102w103w(0) <= wire_altfp_div_pst1_w_datab_range102w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range98w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range108w109w(0) <= wire_altfp_div_pst1_w_datab_range108w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range104w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range114w115w(0) <= wire_altfp_div_pst1_w_datab_range114w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range110w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range120w121w(0) <= wire_altfp_div_pst1_w_datab_range120w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range116w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range126w127w(0) <= wire_altfp_div_pst1_w_datab_range126w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range122w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range132w133w(0) <= wire_altfp_div_pst1_w_datab_range132w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range128w(0);
	wire_altfp_div_pst1_w_lg_w_datab_range138w139w(0) <= wire_altfp_div_pst1_w_datab_range138w(0) OR wire_altfp_div_pst1_w_man_b_not_zero_w_range134w(0);
	a_is_infinity_w <= wire_altfp_div_pst1_w_lg_w_exp_a_all_one_w_range78w222w(0);
	a_is_nan_w <= (exp_a_all_one_w(7) AND man_a_not_zero_w(22));
	a_zero_b_not <= wire_altfp_div_pst1_w_lg_w_exp_b_not_zero_w_range76w256w(0);
	b1_dffe_w <= ( b1_dffe_0);
	b_is_infinity_w <= wire_altfp_div_pst1_w_lg_w_exp_b_all_one_w_range80w224w(0);
	b_is_nan_w <= (exp_b_all_one_w(7) AND man_b_not_zero_w(22));
	bias_addition_overf_w <= wire_bias_addition_overflow;
	bias_addition_w <= wire_bias_addition_result(7 DOWNTO 0);
	both_exp_zeros <= both_exp_zeros_dffe;
	e0_dffe1_wo <= e0_w;
	e0_w <= wire_altsyncram3_q_a;
	e1_w <= ( e1_dffe_1 & e1_dffe_0 & wire_b1_prod_w_lg_w_result_range358w359w);
	exp_a_all_one_w <= ( wire_altfp_div_pst1_w_lg_w_dataa_range71w77w & wire_altfp_div_pst1_w_lg_w_dataa_range61w67w & wire_altfp_div_pst1_w_lg_w_dataa_range51w57w & wire_altfp_div_pst1_w_lg_w_dataa_range41w47w & wire_altfp_div_pst1_w_lg_w_dataa_range31w37w & wire_altfp_div_pst1_w_lg_w_dataa_range21w27w & wire_altfp_div_pst1_w_lg_w_dataa_range11w17w & dataa(23));
	exp_a_not_zero_w <= ( wire_altfp_div_pst1_w_lg_w_dataa_range71w72w & wire_altfp_div_pst1_w_lg_w_dataa_range61w62w & wire_altfp_div_pst1_w_lg_w_dataa_range51w52w & wire_altfp_div_pst1_w_lg_w_dataa_range41w42w & wire_altfp_div_pst1_w_lg_w_dataa_range31w32w & wire_altfp_div_pst1_w_lg_w_dataa_range21w22w & wire_altfp_div_pst1_w_lg_w_dataa_range11w12w & dataa(23));
	exp_add_output_all_one <= ( wire_altfp_div_pst1_w_lg_w_bias_addition_w_range280w297w & wire_altfp_div_pst1_w_lg_w_bias_addition_w_range277w295w & wire_altfp_div_pst1_w_lg_w_bias_addition_w_range274w293w & wire_altfp_div_pst1_w_lg_w_bias_addition_w_range271w291w & wire_altfp_div_pst1_w_lg_w_bias_addition_w_range268w289w & wire_altfp_div_pst1_w_lg_w_bias_addition_w_range265w287w & wire_altfp_div_pst1_w_lg_w_bias_addition_w_range262w285w & bias_addition_w(0));
	exp_add_output_not_zero <= ( wire_altfp_div_pst1_w_lg_w_bias_addition_w_range280w281w & wire_altfp_div_pst1_w_lg_w_bias_addition_w_range277w278w & wire_altfp_div_pst1_w_lg_w_bias_addition_w_range274w275w & wire_altfp_div_pst1_w_lg_w_bias_addition_w_range271w272w & wire_altfp_div_pst1_w_lg_w_bias_addition_w_range268w269w & wire_altfp_div_pst1_w_lg_w_bias_addition_w_range265w266w & wire_altfp_div_pst1_w_lg_w_bias_addition_w_range262w263w & bias_addition_w(0));
	exp_b_all_one_w <= ( wire_altfp_div_pst1_w_lg_w_datab_range74w79w & wire_altfp_div_pst1_w_lg_w_datab_range64w69w & wire_altfp_div_pst1_w_lg_w_datab_range54w59w & wire_altfp_div_pst1_w_lg_w_datab_range44w49w & wire_altfp_div_pst1_w_lg_w_datab_range34w39w & wire_altfp_div_pst1_w_lg_w_datab_range24w29w & wire_altfp_div_pst1_w_lg_w_datab_range14w19w & datab(23));
	exp_b_not_zero_w <= ( wire_altfp_div_pst1_w_lg_w_datab_range74w75w & wire_altfp_div_pst1_w_lg_w_datab_range64w65w & wire_altfp_div_pst1_w_lg_w_datab_range54w55w & wire_altfp_div_pst1_w_lg_w_datab_range44w45w & wire_altfp_div_pst1_w_lg_w_datab_range34w35w & wire_altfp_div_pst1_w_lg_w_datab_range24w25w & wire_altfp_div_pst1_w_lg_w_datab_range14w15w & datab(23));
	exp_result_mux_out <= wire_exp_result_muxa_dataout;
	exp_result_mux_sel_w <= ((((a_zero_b_not_dffe_1 OR b_is_infinity_dffe_1) OR wire_altfp_div_pst1_w_lg_w_lg_bias_addition_overf_w304w312w(0)) OR (((NOT exp_add_output_not_zero(7)) AND wire_altfp_div_pst1_w_lg_bias_addition_overf_w304w(0)) AND wire_altfp_div_pst1_w_lg_exp_sign_w303w(0))) AND wire_nan_pipe_dffe_1_w_lg_q308w(0));
	exp_result_w <= (wire_altfp_div_pst1_w_lg_w_lg_w_lg_bias_addition_overf_w304w305w306w OR wire_altfp_div_pst1_w302w);
	exp_sign_w <= wire_bias_addition_result(8);
	exp_sub_a_w <= ( "0" & dataa(30 DOWNTO 23));
	exp_sub_b_w <= ( "0" & datab(30 DOWNTO 23));
	exp_sub_w <= wire_exp_sub_result;
	frac_a_smaller_dffe1_wi <= frac_a_smaller_w;
	frac_a_smaller_dffe1_wo <= frac_a_smaller_dffe1;
	frac_a_smaller_w <= wire_cmpr2_alb;
	guard_bit <= wire_q_partial_1_result(22);
	man_a_adjusted_w <= wire_man_a_adjusteda_dataout;
	man_a_dffe1_wi <= dataa(22 DOWNTO 0);
	man_a_dffe1_wo <= man_a_dffe1_dffe1;
	man_a_not_zero_w <= ( wire_altfp_div_pst1_w_lg_w_dataa_range213w214w & wire_altfp_div_pst1_w_lg_w_dataa_range207w208w & wire_altfp_div_pst1_w_lg_w_dataa_range201w202w & wire_altfp_div_pst1_w_lg_w_dataa_range195w196w & wire_altfp_div_pst1_w_lg_w_dataa_range189w190w & wire_altfp_div_pst1_w_lg_w_dataa_range183w184w & wire_altfp_div_pst1_w_lg_w_dataa_range177w178w & wire_altfp_div_pst1_w_lg_w_dataa_range171w172w & wire_altfp_div_pst1_w_lg_w_dataa_range165w166w & wire_altfp_div_pst1_w_lg_w_dataa_range159w160w & wire_altfp_div_pst1_w_lg_w_dataa_range153w154w & wire_altfp_div_pst1_w_lg_w_dataa_range147w148w & wire_altfp_div_pst1_w_lg_w_dataa_range141w142w & wire_altfp_div_pst1_w_lg_w_dataa_range135w136w & wire_altfp_div_pst1_w_lg_w_dataa_range129w130w & wire_altfp_div_pst1_w_lg_w_dataa_range123w124w & wire_altfp_div_pst1_w_lg_w_dataa_range117w118w & wire_altfp_div_pst1_w_lg_w_dataa_range111w112w & wire_altfp_div_pst1_w_lg_w_dataa_range105w106w & wire_altfp_div_pst1_w_lg_w_dataa_range99w100w & wire_altfp_div_pst1_w_lg_w_dataa_range93w94w & wire_altfp_div_pst1_w_lg_w_dataa_range87w88w & dataa(0));
	man_b_adjusted_w <= ( "1" & man_b_dffe1_wo);
	man_b_dffe1_wi <= datab(22 DOWNTO 0);
	man_b_dffe1_wo <= man_b_dffe1_dffe1;
	man_b_not_zero_w <= ( wire_altfp_div_pst1_w_lg_w_datab_range216w217w & wire_altfp_div_pst1_w_lg_w_datab_range210w211w & wire_altfp_div_pst1_w_lg_w_datab_range204w205w & wire_altfp_div_pst1_w_lg_w_datab_range198w199w & wire_altfp_div_pst1_w_lg_w_datab_range192w193w & wire_altfp_div_pst1_w_lg_w_datab_range186w187w & wire_altfp_div_pst1_w_lg_w_datab_range180w181w & wire_altfp_div_pst1_w_lg_w_datab_range174w175w & wire_altfp_div_pst1_w_lg_w_datab_range168w169w & wire_altfp_div_pst1_w_lg_w_datab_range162w163w & wire_altfp_div_pst1_w_lg_w_datab_range156w157w & wire_altfp_div_pst1_w_lg_w_datab_range150w151w & wire_altfp_div_pst1_w_lg_w_datab_range144w145w & wire_altfp_div_pst1_w_lg_w_datab_range138w139w & wire_altfp_div_pst1_w_lg_w_datab_range132w133w & wire_altfp_div_pst1_w_lg_w_datab_range126w127w & wire_altfp_div_pst1_w_lg_w_datab_range120w121w & wire_altfp_div_pst1_w_lg_w_datab_range114w115w & wire_altfp_div_pst1_w_lg_w_datab_range108w109w & wire_altfp_div_pst1_w_lg_w_datab_range102w103w & wire_altfp_div_pst1_w_lg_w_datab_range96w97w & wire_altfp_div_pst1_w_lg_w_datab_range90w91w & datab(0));
	man_result_dffe_wi <= man_result_w;
	man_result_dffe_wo <= man_result_dffe;
	man_result_mux_select <= (((((over_under_dffe_2 OR a_zero_b_not_dffe_4) OR nan_pipe_dffe_4) OR b_is_infinity_dffe_4) OR a_is_infinity_dffe_4) OR divbyzero_pipe_dffe_4);
	man_result_w <= wire_man_result_muxa_dataout;
	man_zeros_w <= (OTHERS => '0');
	overflow_ones_w <= (OTHERS => '1');
	overflow_underflow <= (overflow_w OR underflow_w);
	overflow_w <= (wire_altfp_div_pst1_w_lg_bias_addition_overf_w323w(0) AND ((wire_nan_pipe_dffe_1_w_lg_q308w(0) AND wire_a_is_infinity_dffe_1_w_lg_q318w(0)) AND wire_divbyzero_pipe_dffe_1_w_lg_q317w(0)));
	quotient_accumulate_w <= ( quotient_k_dffe_0 & "00000000000000" & quotient_j_dffe & "00000000000000");
	quotient_process_cin_w <= (round_bit AND (guard_bit OR sticky_bits(4)));
	remainder_j_w <= ( wire_remainder_sub_0_result(35 DOWNTO 0) & "00000000000000" & wire_a1_prod_result(34 DOWNTO 0) & "000000000000000");
	result <= ( sign_pipe_dffe_5 & exp_result_dffe_3 & man_result_dffe_wo);
	round_bit <= wire_q_partial_1_result(21);
	select_bias_out_2_w <= wire_select_bias_2a_dataout;
	select_bias_out_w <= wire_select_biasa_dataout;
	sticky_bits <= ( wire_q_partial_1_w_lg_w_result_range416w417w & wire_q_partial_1_w_lg_w_result_range413w414w & wire_q_partial_1_w_lg_w_result_range410w411w & wire_q_partial_1_w_lg_w_result_range407w408w & wire_q_partial_1_result(16));
	underflow_w <= ((((wire_altfp_div_pst1_w_lg_w_lg_bias_addition_overf_w304w312w(0) OR (((NOT exp_add_output_not_zero(7)) AND wire_altfp_div_pst1_w_lg_bias_addition_overf_w304w(0)) AND wire_altfp_div_pst1_w_lg_exp_sign_w303w(0))) AND wire_nan_pipe_dffe_1_w_lg_q308w(0)) AND wire_a_zero_b_not_dffe_1_w_lg_q326w(0)) AND wire_b_is_infinity_dffe_1_w_lg_q325w(0));
	underflow_zeros_w <= (OTHERS => '0');
	value_add_one_w <= "001111111";
	value_normal_w <= "001111110";
	value_zero_w <= (OTHERS => '0');
	wire_altfp_div_pst1_w_bias_addition_w_range262w(0) <= bias_addition_w(1);
	wire_altfp_div_pst1_w_bias_addition_w_range265w(0) <= bias_addition_w(2);
	wire_altfp_div_pst1_w_bias_addition_w_range268w(0) <= bias_addition_w(3);
	wire_altfp_div_pst1_w_bias_addition_w_range271w(0) <= bias_addition_w(4);
	wire_altfp_div_pst1_w_bias_addition_w_range274w(0) <= bias_addition_w(5);
	wire_altfp_div_pst1_w_bias_addition_w_range277w(0) <= bias_addition_w(6);
	wire_altfp_div_pst1_w_bias_addition_w_range280w(0) <= bias_addition_w(7);
	wire_altfp_div_pst1_w_dataa_range141w(0) <= dataa(10);
	wire_altfp_div_pst1_w_dataa_range147w(0) <= dataa(11);
	wire_altfp_div_pst1_w_dataa_range153w(0) <= dataa(12);
	wire_altfp_div_pst1_w_dataa_range159w(0) <= dataa(13);
	wire_altfp_div_pst1_w_dataa_range165w(0) <= dataa(14);
	wire_altfp_div_pst1_w_dataa_range171w(0) <= dataa(15);
	wire_altfp_div_pst1_w_dataa_range177w(0) <= dataa(16);
	wire_altfp_div_pst1_w_dataa_range183w(0) <= dataa(17);
	wire_altfp_div_pst1_w_dataa_range189w(0) <= dataa(18);
	wire_altfp_div_pst1_w_dataa_range195w(0) <= dataa(19);
	wire_altfp_div_pst1_w_dataa_range87w(0) <= dataa(1);
	wire_altfp_div_pst1_w_dataa_range201w(0) <= dataa(20);
	wire_altfp_div_pst1_w_dataa_range207w(0) <= dataa(21);
	wire_altfp_div_pst1_w_dataa_range213w(0) <= dataa(22);
	wire_altfp_div_pst1_w_dataa_range11w(0) <= dataa(24);
	wire_altfp_div_pst1_w_dataa_range21w(0) <= dataa(25);
	wire_altfp_div_pst1_w_dataa_range31w(0) <= dataa(26);
	wire_altfp_div_pst1_w_dataa_range41w(0) <= dataa(27);
	wire_altfp_div_pst1_w_dataa_range51w(0) <= dataa(28);
	wire_altfp_div_pst1_w_dataa_range61w(0) <= dataa(29);
	wire_altfp_div_pst1_w_dataa_range93w(0) <= dataa(2);
	wire_altfp_div_pst1_w_dataa_range71w(0) <= dataa(30);
	wire_altfp_div_pst1_w_dataa_range99w(0) <= dataa(3);
	wire_altfp_div_pst1_w_dataa_range105w(0) <= dataa(4);
	wire_altfp_div_pst1_w_dataa_range111w(0) <= dataa(5);
	wire_altfp_div_pst1_w_dataa_range117w(0) <= dataa(6);
	wire_altfp_div_pst1_w_dataa_range123w(0) <= dataa(7);
	wire_altfp_div_pst1_w_dataa_range129w(0) <= dataa(8);
	wire_altfp_div_pst1_w_dataa_range135w(0) <= dataa(9);
	wire_altfp_div_pst1_w_datab_range144w(0) <= datab(10);
	wire_altfp_div_pst1_w_datab_range150w(0) <= datab(11);
	wire_altfp_div_pst1_w_datab_range156w(0) <= datab(12);
	wire_altfp_div_pst1_w_datab_range162w(0) <= datab(13);
	wire_altfp_div_pst1_w_datab_range168w(0) <= datab(14);
	wire_altfp_div_pst1_w_datab_range174w(0) <= datab(15);
	wire_altfp_div_pst1_w_datab_range180w(0) <= datab(16);
	wire_altfp_div_pst1_w_datab_range186w(0) <= datab(17);
	wire_altfp_div_pst1_w_datab_range192w(0) <= datab(18);
	wire_altfp_div_pst1_w_datab_range198w(0) <= datab(19);
	wire_altfp_div_pst1_w_datab_range90w(0) <= datab(1);
	wire_altfp_div_pst1_w_datab_range204w(0) <= datab(20);
	wire_altfp_div_pst1_w_datab_range210w(0) <= datab(21);
	wire_altfp_div_pst1_w_datab_range216w(0) <= datab(22);
	wire_altfp_div_pst1_w_datab_range14w(0) <= datab(24);
	wire_altfp_div_pst1_w_datab_range24w(0) <= datab(25);
	wire_altfp_div_pst1_w_datab_range34w(0) <= datab(26);
	wire_altfp_div_pst1_w_datab_range44w(0) <= datab(27);
	wire_altfp_div_pst1_w_datab_range54w(0) <= datab(28);
	wire_altfp_div_pst1_w_datab_range64w(0) <= datab(29);
	wire_altfp_div_pst1_w_datab_range96w(0) <= datab(2);
	wire_altfp_div_pst1_w_datab_range74w(0) <= datab(30);
	wire_altfp_div_pst1_w_datab_range102w(0) <= datab(3);
	wire_altfp_div_pst1_w_datab_range108w(0) <= datab(4);
	wire_altfp_div_pst1_w_datab_range114w(0) <= datab(5);
	wire_altfp_div_pst1_w_datab_range120w(0) <= datab(6);
	wire_altfp_div_pst1_w_datab_range126w(0) <= datab(7);
	wire_altfp_div_pst1_w_datab_range132w(0) <= datab(8);
	wire_altfp_div_pst1_w_datab_range138w(0) <= datab(9);
	wire_altfp_div_pst1_w_e1_w_range360w <= e1_w(16 DOWNTO 0);
	wire_altfp_div_pst1_w_e1_w_range368w <= e1_w(33 DOWNTO 17);
	wire_altfp_div_pst1_w_exp_a_all_one_w_range7w(0) <= exp_a_all_one_w(0);
	wire_altfp_div_pst1_w_exp_a_all_one_w_range18w(0) <= exp_a_all_one_w(1);
	wire_altfp_div_pst1_w_exp_a_all_one_w_range28w(0) <= exp_a_all_one_w(2);
	wire_altfp_div_pst1_w_exp_a_all_one_w_range38w(0) <= exp_a_all_one_w(3);
	wire_altfp_div_pst1_w_exp_a_all_one_w_range48w(0) <= exp_a_all_one_w(4);
	wire_altfp_div_pst1_w_exp_a_all_one_w_range58w(0) <= exp_a_all_one_w(5);
	wire_altfp_div_pst1_w_exp_a_all_one_w_range68w(0) <= exp_a_all_one_w(6);
	wire_altfp_div_pst1_w_exp_a_all_one_w_range78w(0) <= exp_a_all_one_w(7);
	wire_altfp_div_pst1_w_exp_a_not_zero_w_range2w(0) <= exp_a_not_zero_w(0);
	wire_altfp_div_pst1_w_exp_a_not_zero_w_range13w(0) <= exp_a_not_zero_w(1);
	wire_altfp_div_pst1_w_exp_a_not_zero_w_range23w(0) <= exp_a_not_zero_w(2);
	wire_altfp_div_pst1_w_exp_a_not_zero_w_range33w(0) <= exp_a_not_zero_w(3);
	wire_altfp_div_pst1_w_exp_a_not_zero_w_range43w(0) <= exp_a_not_zero_w(4);
	wire_altfp_div_pst1_w_exp_a_not_zero_w_range53w(0) <= exp_a_not_zero_w(5);
	wire_altfp_div_pst1_w_exp_a_not_zero_w_range63w(0) <= exp_a_not_zero_w(6);
	wire_altfp_div_pst1_w_exp_a_not_zero_w_range73w(0) <= exp_a_not_zero_w(7);
	wire_altfp_div_pst1_w_exp_add_output_all_one_range283w(0) <= exp_add_output_all_one(0);
	wire_altfp_div_pst1_w_exp_add_output_all_one_range286w(0) <= exp_add_output_all_one(1);
	wire_altfp_div_pst1_w_exp_add_output_all_one_range288w(0) <= exp_add_output_all_one(2);
	wire_altfp_div_pst1_w_exp_add_output_all_one_range290w(0) <= exp_add_output_all_one(3);
	wire_altfp_div_pst1_w_exp_add_output_all_one_range292w(0) <= exp_add_output_all_one(4);
	wire_altfp_div_pst1_w_exp_add_output_all_one_range294w(0) <= exp_add_output_all_one(5);
	wire_altfp_div_pst1_w_exp_add_output_all_one_range296w(0) <= exp_add_output_all_one(6);
	wire_altfp_div_pst1_w_exp_add_output_all_one_range298w(0) <= exp_add_output_all_one(7);
	wire_altfp_div_pst1_w_exp_add_output_not_zero_range260w(0) <= exp_add_output_not_zero(0);
	wire_altfp_div_pst1_w_exp_add_output_not_zero_range264w(0) <= exp_add_output_not_zero(1);
	wire_altfp_div_pst1_w_exp_add_output_not_zero_range267w(0) <= exp_add_output_not_zero(2);
	wire_altfp_div_pst1_w_exp_add_output_not_zero_range270w(0) <= exp_add_output_not_zero(3);
	wire_altfp_div_pst1_w_exp_add_output_not_zero_range273w(0) <= exp_add_output_not_zero(4);
	wire_altfp_div_pst1_w_exp_add_output_not_zero_range276w(0) <= exp_add_output_not_zero(5);
	wire_altfp_div_pst1_w_exp_add_output_not_zero_range279w(0) <= exp_add_output_not_zero(6);
	wire_altfp_div_pst1_w_exp_b_all_one_w_range9w(0) <= exp_b_all_one_w(0);
	wire_altfp_div_pst1_w_exp_b_all_one_w_range20w(0) <= exp_b_all_one_w(1);
	wire_altfp_div_pst1_w_exp_b_all_one_w_range30w(0) <= exp_b_all_one_w(2);
	wire_altfp_div_pst1_w_exp_b_all_one_w_range40w(0) <= exp_b_all_one_w(3);
	wire_altfp_div_pst1_w_exp_b_all_one_w_range50w(0) <= exp_b_all_one_w(4);
	wire_altfp_div_pst1_w_exp_b_all_one_w_range60w(0) <= exp_b_all_one_w(5);
	wire_altfp_div_pst1_w_exp_b_all_one_w_range70w(0) <= exp_b_all_one_w(6);
	wire_altfp_div_pst1_w_exp_b_all_one_w_range80w(0) <= exp_b_all_one_w(7);
	wire_altfp_div_pst1_w_exp_b_not_zero_w_range5w(0) <= exp_b_not_zero_w(0);
	wire_altfp_div_pst1_w_exp_b_not_zero_w_range16w(0) <= exp_b_not_zero_w(1);
	wire_altfp_div_pst1_w_exp_b_not_zero_w_range26w(0) <= exp_b_not_zero_w(2);
	wire_altfp_div_pst1_w_exp_b_not_zero_w_range36w(0) <= exp_b_not_zero_w(3);
	wire_altfp_div_pst1_w_exp_b_not_zero_w_range46w(0) <= exp_b_not_zero_w(4);
	wire_altfp_div_pst1_w_exp_b_not_zero_w_range56w(0) <= exp_b_not_zero_w(5);
	wire_altfp_div_pst1_w_exp_b_not_zero_w_range66w(0) <= exp_b_not_zero_w(6);
	wire_altfp_div_pst1_w_exp_b_not_zero_w_range76w(0) <= exp_b_not_zero_w(7);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range82w(0) <= man_a_not_zero_w(0);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range143w(0) <= man_a_not_zero_w(10);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range149w(0) <= man_a_not_zero_w(11);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range155w(0) <= man_a_not_zero_w(12);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range161w(0) <= man_a_not_zero_w(13);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range167w(0) <= man_a_not_zero_w(14);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range173w(0) <= man_a_not_zero_w(15);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range179w(0) <= man_a_not_zero_w(16);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range185w(0) <= man_a_not_zero_w(17);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range191w(0) <= man_a_not_zero_w(18);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range197w(0) <= man_a_not_zero_w(19);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range89w(0) <= man_a_not_zero_w(1);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range203w(0) <= man_a_not_zero_w(20);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range209w(0) <= man_a_not_zero_w(21);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range215w(0) <= man_a_not_zero_w(22);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range95w(0) <= man_a_not_zero_w(2);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range101w(0) <= man_a_not_zero_w(3);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range107w(0) <= man_a_not_zero_w(4);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range113w(0) <= man_a_not_zero_w(5);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range119w(0) <= man_a_not_zero_w(6);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range125w(0) <= man_a_not_zero_w(7);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range131w(0) <= man_a_not_zero_w(8);
	wire_altfp_div_pst1_w_man_a_not_zero_w_range137w(0) <= man_a_not_zero_w(9);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range85w(0) <= man_b_not_zero_w(0);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range146w(0) <= man_b_not_zero_w(10);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range152w(0) <= man_b_not_zero_w(11);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range158w(0) <= man_b_not_zero_w(12);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range164w(0) <= man_b_not_zero_w(13);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range170w(0) <= man_b_not_zero_w(14);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range176w(0) <= man_b_not_zero_w(15);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range182w(0) <= man_b_not_zero_w(16);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range188w(0) <= man_b_not_zero_w(17);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range194w(0) <= man_b_not_zero_w(18);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range200w(0) <= man_b_not_zero_w(19);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range92w(0) <= man_b_not_zero_w(1);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range206w(0) <= man_b_not_zero_w(20);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range212w(0) <= man_b_not_zero_w(21);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range218w(0) <= man_b_not_zero_w(22);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range98w(0) <= man_b_not_zero_w(2);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range104w(0) <= man_b_not_zero_w(3);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range110w(0) <= man_b_not_zero_w(4);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range116w(0) <= man_b_not_zero_w(5);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range122w(0) <= man_b_not_zero_w(6);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range128w(0) <= man_b_not_zero_w(7);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range134w(0) <= man_b_not_zero_w(8);
	wire_altfp_div_pst1_w_man_b_not_zero_w_range140w(0) <= man_b_not_zero_w(9);
	wire_altfp_div_pst1_w_remainder_j_w_range363w <= remainder_j_w(49 DOWNTO 0);
	wire_altfp_div_pst1_w_sticky_bits_range405w(0) <= sticky_bits(0);
	wire_altfp_div_pst1_w_sticky_bits_range409w(0) <= sticky_bits(1);
	wire_altfp_div_pst1_w_sticky_bits_range412w(0) <= sticky_bits(2);
	wire_altfp_div_pst1_w_sticky_bits_range415w(0) <= sticky_bits(3);
	wire_altfp_div_pst1_w_w_quotient_accumulate_w_range385w_range386w <= quotient_accumulate_w(30 DOWNTO 14);
	altsyncram3 :  altsyncram
	  GENERIC MAP (
		INIT_FILE => "alt_float_div.hex",
		OPERATION_MODE => "ROM",
		WIDTH_A => 9,
		WIDTHAD_A => 9,
		INTENDED_DEVICE_FAMILY => "Cyclone V"
	  )
	  PORT MAP ( 
		address_a => datab(22 DOWNTO 14),
		clock0 => clock,
		clocken0 => clk_en,
		q_a => wire_altsyncram3_q_a
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN a_is_infinity_dffe_0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN a_is_infinity_dffe_0 <= a_is_infinity_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN a_is_infinity_dffe_1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN a_is_infinity_dffe_1 <= a_is_infinity_dffe_0;
			END IF;
		END IF;
	END PROCESS;
	wire_a_is_infinity_dffe_1_w_lg_q318w(0) <= NOT a_is_infinity_dffe_1;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN a_is_infinity_dffe_2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN a_is_infinity_dffe_2 <= a_is_infinity_dffe_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN a_is_infinity_dffe_3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN a_is_infinity_dffe_3 <= a_is_infinity_dffe_2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN a_is_infinity_dffe_4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN a_is_infinity_dffe_4 <= a_is_infinity_dffe_3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN a_zero_b_not_dffe_0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN a_zero_b_not_dffe_0 <= a_zero_b_not;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN a_zero_b_not_dffe_1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN a_zero_b_not_dffe_1 <= a_zero_b_not_dffe_0;
			END IF;
		END IF;
	END PROCESS;
	wire_a_zero_b_not_dffe_1_w_lg_q326w(0) <= NOT a_zero_b_not_dffe_1;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN a_zero_b_not_dffe_2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN a_zero_b_not_dffe_2 <= a_zero_b_not_dffe_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN a_zero_b_not_dffe_3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN a_zero_b_not_dffe_3 <= a_zero_b_not_dffe_2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN a_zero_b_not_dffe_4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN a_zero_b_not_dffe_4 <= a_zero_b_not_dffe_3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN b1_dffe_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN b1_dffe_0 <= wire_b1_prod_result;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN b_is_infinity_dffe_0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN b_is_infinity_dffe_0 <= b_is_infinity_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN b_is_infinity_dffe_1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN b_is_infinity_dffe_1 <= b_is_infinity_dffe_0;
			END IF;
		END IF;
	END PROCESS;
	wire_b_is_infinity_dffe_1_w_lg_q325w(0) <= NOT b_is_infinity_dffe_1;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN b_is_infinity_dffe_2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN b_is_infinity_dffe_2 <= b_is_infinity_dffe_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN b_is_infinity_dffe_3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN b_is_infinity_dffe_3 <= b_is_infinity_dffe_2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN b_is_infinity_dffe_4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN b_is_infinity_dffe_4 <= b_is_infinity_dffe_3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN both_exp_zeros_dffe <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN both_exp_zeros_dffe <= ((NOT exp_b_not_zero_w(7)) AND wire_altfp_div_pst1_w_lg_w_exp_a_not_zero_w_range73w227w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN divbyzero_pipe_dffe_0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN divbyzero_pipe_dffe_0 <= ((((NOT exp_b_not_zero_w(7)) AND wire_altfp_div_pst1_w_lg_a_is_nan_w234w(0)) AND exp_a_not_zero_w(7)) AND wire_altfp_div_pst1_w_lg_a_is_infinity_w233w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN divbyzero_pipe_dffe_1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN divbyzero_pipe_dffe_1 <= divbyzero_pipe_dffe_0;
			END IF;
		END IF;
	END PROCESS;
	wire_divbyzero_pipe_dffe_1_w_lg_q317w(0) <= NOT divbyzero_pipe_dffe_1;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN divbyzero_pipe_dffe_2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN divbyzero_pipe_dffe_2 <= divbyzero_pipe_dffe_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN divbyzero_pipe_dffe_3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN divbyzero_pipe_dffe_3 <= divbyzero_pipe_dffe_2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN divbyzero_pipe_dffe_4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN divbyzero_pipe_dffe_4 <= divbyzero_pipe_dffe_3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN e1_dffe_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN e1_dffe_0 <= wire_altfp_div_pst1_w_e1_w_range360w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN e1_dffe_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN e1_dffe_1 <= wire_altfp_div_pst1_w_e1_w_range368w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_result_dffe_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_result_dffe_0 <= exp_result_mux_out;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_result_dffe_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_result_dffe_1 <= exp_result_dffe_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_result_dffe_2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_result_dffe_2 <= exp_result_dffe_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_result_dffe_3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_result_dffe_3 <= exp_result_dffe_2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN frac_a_smaller_dffe1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN frac_a_smaller_dffe1 <= frac_a_smaller_dffe1_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_a_dffe1_dffe1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_a_dffe1_dffe1 <= man_a_dffe1_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_b_dffe1_dffe1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_b_dffe1_dffe1 <= man_b_dffe1_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_result_dffe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_result_dffe <= man_result_dffe_wi;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_pipe_dffe_0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_pipe_dffe_0 <= (((a_is_nan_w OR b_is_nan_w) OR (a_is_infinity_w AND b_is_infinity_w)) OR (wire_altfp_div_pst1_w_lg_w_exp_a_not_zero_w_range73w227w(0) AND (NOT exp_b_not_zero_w(7))));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_pipe_dffe_1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_pipe_dffe_1 <= nan_pipe_dffe_0;
			END IF;
		END IF;
	END PROCESS;
	wire_nan_pipe_dffe_1_w_lg_q308w(0) <= NOT nan_pipe_dffe_1;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_pipe_dffe_2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_pipe_dffe_2 <= nan_pipe_dffe_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_pipe_dffe_3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_pipe_dffe_3 <= nan_pipe_dffe_2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_pipe_dffe_4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_pipe_dffe_4 <= nan_pipe_dffe_3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN over_under_dffe_0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN over_under_dffe_0 <= overflow_underflow;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN over_under_dffe_1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN over_under_dffe_1 <= over_under_dffe_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN over_under_dffe_2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN over_under_dffe_2 <= over_under_dffe_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN quotient_j_dffe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN quotient_j_dffe <= wire_q_partial_0_w_result_range373w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN quotient_k_dffe_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN quotient_k_dffe_0 <= wire_altfp_div_pst1_w_w_quotient_accumulate_w_range385w_range386w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN remainder_j_dffe_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN remainder_j_dffe_0 <= wire_altfp_div_pst1_w_remainder_j_w_range363w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN remainder_j_dffe_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN remainder_j_dffe_1 <= remainder_j_dffe_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_pipe_dffe_0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_pipe_dffe_0 <= (dataa(31) XOR datab(31));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_pipe_dffe_1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_pipe_dffe_1 <= sign_pipe_dffe_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_pipe_dffe_2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_pipe_dffe_2 <= sign_pipe_dffe_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_pipe_dffe_3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_pipe_dffe_3 <= sign_pipe_dffe_2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_pipe_dffe_4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_pipe_dffe_4 <= sign_pipe_dffe_3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_pipe_dffe_5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_pipe_dffe_5 <= sign_pipe_dffe_4;
			END IF;
		END IF;
	END PROCESS;
	bias_addition :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => exp_sub_w,
		datab => select_bias_out_2_w,
		overflow => wire_bias_addition_overflow,
		result => wire_bias_addition_result
	  );
	exp_sub :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => exp_sub_a_w,
		datab => exp_sub_b_w,
		result => wire_exp_sub_result
	  );
	wire_quotient_process_dataa <= ( quotient_accumulate_w(61 DOWNTO 45) & "00000000000000");
	wire_quotient_process_datab <= ( "00000000000000" & wire_q_partial_1_result(32 DOWNTO 22) & "111111");
	wire_quotient_process_w_result_range425w <= wire_quotient_process_result(28 DOWNTO 6);
	quotient_process :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 31
	  )
	  PORT MAP ( 
		cin => quotient_process_cin_w,
		dataa => wire_quotient_process_dataa,
		datab => wire_quotient_process_datab,
		result => wire_quotient_process_result
	  );
	wire_remainder_sub_0_dataa <= ( remainder_j_dffe_1(49 DOWNTO 15) & "000000000000000");
	remainder_sub_0 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 50
	  )
	  PORT MAP ( 
		dataa => wire_remainder_sub_0_dataa,
		datab => wire_remainder_mult_0_result(49 DOWNTO 0),
		result => wire_remainder_sub_0_result
	  );
	cmpr2 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 23
	  )
	  PORT MAP ( 
		alb => wire_cmpr2_alb,
		dataa => dataa(22 DOWNTO 0),
		datab => datab(22 DOWNTO 0)
	  );
	wire_a1_prod_datab <= ( "1" & e0_dffe1_wo);
	a1_prod :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 25,
		LPM_WIDTHB => 10,
		LPM_WIDTHP => 35,
		lpm_hint => "DEDICATED_MULTIPLIER_CIRCUITRY=YES"
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => man_a_adjusted_w,
		datab => wire_a1_prod_datab,
		result => wire_a1_prod_result
	  );
	loop2 : FOR i IN 0 TO 16 GENERATE 
		wire_b1_prod_w_lg_w_result_range358w359w(i) <= NOT wire_b1_prod_w_result_range358w(i);
	END GENERATE loop2;
	wire_b1_prod_datab <= ( "1" & e0_dffe1_wo);
	wire_b1_prod_w_result_range358w <= wire_b1_prod_result(33 DOWNTO 17);
	b1_prod :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 24,
		LPM_WIDTHB => 10,
		LPM_WIDTHP => 34,
		lpm_hint => "DEDICATED_MULTIPLIER_CIRCUITRY=YES"
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => man_b_adjusted_w,
		datab => wire_b1_prod_datab,
		result => wire_b1_prod_result
	  );
	wire_q_partial_0_w_result_range373w <= wire_q_partial_0_result(32 DOWNTO 16);
	q_partial_0 :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 17,
		LPM_WIDTHB => 17,
		LPM_WIDTHP => 34,
		lpm_hint => "DEDICATED_MULTIPLIER_CIRCUITRY=YES"
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => remainder_j_w(49 DOWNTO 33),
		datab => e1_w(16 DOWNTO 0),
		result => wire_q_partial_0_result
	  );
	wire_q_partial_1_w_lg_w_result_range407w408w(0) <= wire_q_partial_1_w_result_range407w(0) OR wire_altfp_div_pst1_w_sticky_bits_range405w(0);
	wire_q_partial_1_w_lg_w_result_range410w411w(0) <= wire_q_partial_1_w_result_range410w(0) OR wire_altfp_div_pst1_w_sticky_bits_range409w(0);
	wire_q_partial_1_w_lg_w_result_range413w414w(0) <= wire_q_partial_1_w_result_range413w(0) OR wire_altfp_div_pst1_w_sticky_bits_range412w(0);
	wire_q_partial_1_w_lg_w_result_range416w417w(0) <= wire_q_partial_1_w_result_range416w(0) OR wire_altfp_div_pst1_w_sticky_bits_range415w(0);
	wire_q_partial_1_w_result_range407w(0) <= wire_q_partial_1_result(17);
	wire_q_partial_1_w_result_range410w(0) <= wire_q_partial_1_result(18);
	wire_q_partial_1_w_result_range413w(0) <= wire_q_partial_1_result(19);
	wire_q_partial_1_w_result_range416w(0) <= wire_q_partial_1_result(20);
	q_partial_1 :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 17,
		LPM_WIDTHB => 17,
		LPM_WIDTHP => 34,
		lpm_hint => "DEDICATED_MULTIPLIER_CIRCUITRY=YES"
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => remainder_j_w(99 DOWNTO 83),
		datab => e1_w(50 DOWNTO 34),
		result => wire_q_partial_1_result
	  );
	remainder_mult_0 :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 34,
		LPM_WIDTHB => 17,
		LPM_WIDTHP => 51,
		lpm_hint => "DEDICATED_MULTIPLIER_CIRCUITRY=YES"
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => b1_dffe_w(33 DOWNTO 0),
		datab => wire_q_partial_0_result(32 DOWNTO 16),
		result => wire_remainder_mult_0_result
	  );
	wire_exp_result_muxa_dataout <= underflow_zeros_w WHEN exp_result_mux_sel_w = '1'  ELSE exp_result_w;
	wire_man_a_adjusteda_dataout <= ( "1" & man_a_dffe1_wo & "0") WHEN frac_a_smaller_dffe1_wo = '1'  ELSE ( "0" & "1" & man_a_dffe1_wo);
	wire_man_result_muxa_dataout <= ( nan_pipe_dffe_4 & man_zeros_w(21 DOWNTO 0)) WHEN man_result_mux_select = '1'  ELSE wire_quotient_process_result(28 DOWNTO 6);
	wire_select_bias_2a_dataout <= value_zero_w WHEN both_exp_zeros = '1'  ELSE select_bias_out_w;
	wire_select_biasa_dataout <= value_normal_w WHEN frac_a_smaller_dffe1_wo = '1'  ELSE value_add_one_w;

 END RTL; --alt_float_div_altfp_div_pst_jcf

--synthesis_resources = altsyncram 1 lpm_add_sub 4 lpm_compare 1 lpm_mult 5 mux21 74 reg 339 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  alt_float_div_altfp_div_i3i IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clk_en	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC;
		 dataa	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 datab	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0)
	 ); 
 END alt_float_div_altfp_div_i3i;

 ARCHITECTURE RTL OF alt_float_div_altfp_div_i3i IS

	 SIGNAL  wire_altfp_div_pst1_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 COMPONENT  alt_float_div_altfp_div_pst_jcf
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clk_en	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC;
		dataa	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		datab	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		result	:	OUT  STD_LOGIC_VECTOR(31 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	result <= wire_altfp_div_pst1_result;
	altfp_div_pst1 :  alt_float_div_altfp_div_pst_jcf
	  PORT MAP ( 
		aclr => aclr,
		clk_en => clk_en,
		clock => clock,
		dataa => dataa,
		datab => datab,
		result => wire_altfp_div_pst1_result
	  );

 END RTL; --alt_float_div_altfp_div_i3i
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY alt_float_div IS
	PORT
	(
		aclr		: IN STD_LOGIC ;
		clk_en		: IN STD_LOGIC ;
		clock		: IN STD_LOGIC ;
		dataa		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		datab		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END alt_float_div;


ARCHITECTURE RTL OF alt_float_div IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (31 DOWNTO 0);



	COMPONENT alt_float_div_altfp_div_i3i
	PORT (
			aclr	: IN STD_LOGIC ;
			clk_en	: IN STD_LOGIC ;
			clock	: IN STD_LOGIC ;
			dataa	: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			datab	: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			result	: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	result    <= sub_wire0(31 DOWNTO 0);

	alt_float_div_altfp_div_i3i_component : alt_float_div_altfp_div_i3i
	PORT MAP (
		aclr => aclr,
		clk_en => clk_en,
		clock => clock,
		dataa => dataa,
		datab => datab,
		result => sub_wire0
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: DENORMAL_SUPPORT STRING "NO"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: CONSTANT: OPTIMIZE STRING "AREA"
-- Retrieval info: CONSTANT: PIPELINE NUMERIC "6"
-- Retrieval info: CONSTANT: REDUCED_FUNCTIONALITY STRING "NO"
-- Retrieval info: CONSTANT: WIDTH_EXP NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_MAN NUMERIC "23"
-- Retrieval info: USED_PORT: aclr 0 0 0 0 INPUT NODEFVAL "aclr"
-- Retrieval info: USED_PORT: clk_en 0 0 0 0 INPUT NODEFVAL "clk_en"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: USED_PORT: dataa 0 0 32 0 INPUT NODEFVAL "dataa[31..0]"
-- Retrieval info: USED_PORT: datab 0 0 32 0 INPUT NODEFVAL "datab[31..0]"
-- Retrieval info: USED_PORT: result 0 0 32 0 OUTPUT NODEFVAL "result[31..0]"
-- Retrieval info: CONNECT: @aclr 0 0 0 0 aclr 0 0 0 0
-- Retrieval info: CONNECT: @clk_en 0 0 0 0 clk_en 0 0 0 0
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: CONNECT: @dataa 0 0 32 0 dataa 0 0 32 0
-- Retrieval info: CONNECT: @datab 0 0 32 0 datab 0 0 32 0
-- Retrieval info: CONNECT: result 0 0 32 0 @result 0 0 32 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL alt_float_div.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL alt_float_div.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL alt_float_div.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL alt_float_div.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL alt_float_div_inst.vhd FALSE
