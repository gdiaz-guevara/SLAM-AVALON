-- altera vhdl_input_version vhdl_2008
------------------------------------------------
LIBRARY ieee;
	USE ieee.std_logic_1164.all;
	USE ieee.numeric_std.all;

------------------------------------------------
PACKAGE my_package IS
	--===================================================
	--             CONSTANT DECLARATIONS
	--===================================================
	CONSTANT DATA_WIDTH					:	INTEGER																:=	32;
	CONSTANT ADDR_AVALON_WIDTH			:	INTEGER																:=	15; --7;
	--CONSTANT ADDR_WIDTH					:	INTEGER															:=	4; 
	CONSTANT IPMEM_DATA_WIDTH			:	INTEGER																:=	108; 
		
	CONSTANT INPUT_DATA_ADDR_WIDTH	:	INTEGER																:=	14; --4;
	CONSTANT QUADRANT_ADDR_WIDTH		:	INTEGER																:=	11; --4;
	CONSTANT VOXEL_ADDR_WIDTH			:	INTEGER																:=	8;  --3;
	CONSTANT MAP_ADDR_WIDTH				:	INTEGER																:=	13;--4;
	
--	CONSTANT ADDR_WIDTH				:	INTEGER																:=	15; -- 15 para prueba grande
--	CONSTANT ADDR_AVALON_WIDTH		:	INTEGER																:=	18;  -- 18 para prueba grande
	
	CONSTANT LATENCY_WIDTH			:	INTEGER																:=	8;
	
	CONSTANT	ZEROS							:	STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0) 					:= (OTHERS => '0');
	CONSTANT	ONE_BIN						:	STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0) 					:= "00000000000000000000000000000001";	
	CONSTANT	ONE_HUNDRED_BIN			:	STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0) 					:= "00000000000000000000000001100100";
	CONSTANT	FP_THOUSAND					:	STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0)					:= "01000100011110100000000000000000"; -- 1000.00
	CONSTANT Z_THRESHOLD					:	STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0) 					:= "11111111111111111111111010000100"; -- 0d-380°
	CONSTANT X_MAP_THRESHOLD			:	STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0) 					:= "00111101100001010001111010111000";	-- 0.065
	CONSTANT Y_MAP_THRESHOLD			:	STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0) 					:= "00111101100001010001111010111000";	-- 0.065
	CONSTANT Z_MAP_THRESHOLD			:	STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0) 					:= "00111101100001010001111010111000";	-- 0.065
	
	CONSTANT	MINUS_ONE_BIN				:	STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0) 					:= (OTHERS => '1'); -- -1
	CONSTANT FLOAT_MULT_LATENCY		:	UNSIGNED(LATENCY_WIDTH-1 DOWNTO 0)		 					:= to_unsigned(5,LATENCY_WIDTH); -- 5
	CONSTANT FLOAT_DIV_LATENCY			:	UNSIGNED(LATENCY_WIDTH-1 DOWNTO 0)		 					:= to_unsigned(6,LATENCY_WIDTH); -- 6
	CONSTANT FLOAT_ADD_LATENCY			:	UNSIGNED(LATENCY_WIDTH-1 DOWNTO 0)		 					:= to_unsigned(7,LATENCY_WIDTH); -- 7
	CONSTANT FLOAT2INT_LATENCY			:	UNSIGNED(LATENCY_WIDTH-1 DOWNTO 0)							:= to_unsigned(6,LATENCY_WIDTH); -- 6
	CONSTANT FLOAT_COMP_LATENCY		:	UNSIGNED(LATENCY_WIDTH-1 DOWNTO 0)							:= to_unsigned(3,LATENCY_WIDTH); -- 3
	--CONSTANT	PADDING_Z_ADDR2DATA_UN	:	UNSIGNED((DATA_WIDTH-ADDR_WIDTH)-1 DOWNTO 0)			 	:= (OTHERS => '0');	
	--CONSTANT	PADDING_Z_ADDR2DATA		:	STD_LOGIC_VECTOR((DATA_WIDTH-ADDR_WIDTH)-1 DOWNTO 0)	:= (OTHERS => '0');	
	CONSTANT	PADDING_Z_ADDRQ2DATA		:	STD_LOGIC_VECTOR((DATA_WIDTH-QUADRANT_ADDR_WIDTH)-1 DOWNTO 0)	:= (OTHERS => '0');	
	CONSTANT	PADDING_Z_MAP_ADDR2DATA	:	STD_LOGIC_VECTOR((DATA_WIDTH-MAP_ADDR_WIDTH)-1 DOWNTO 0)	:= (OTHERS => '0');	
	CONSTANT	PADDING_Z_ADDRQ2DATA_UN	:	UNSIGNED((DATA_WIDTH-QUADRANT_ADDR_WIDTH)-1 DOWNTO 0)	:= (OTHERS => '0');	
	CONSTANT PADDING_BIT					:	STD_LOGIC_VECTOR(DATA_WIDTH-2 DOWNTO 0)					:= (OTHERS => '0');
	CONSTANT PADDING_WORD				:	STD_LOGIC_VECTOR(95 DOWNTO 0)									:= (OTHERS => '0');
	CONSTANT	PADDING_AV2ARRAY_UNSIGNED:	UNSIGNED((ADDR_AVALON_WIDTH-INPUT_DATA_ADDR_WIDTH)-1 DOWNTO 0)	:= (OTHERS => '0');	
	CONSTANT	PADDING_POINT2_IPMEM		:	STD_LOGIC_VECTOR(11 DOWNTO 0)							:= (OTHERS => '0');	
	CONSTANT	MAX_VOXEL_SIZE				:	STD_LOGIC_VECTOR(VOXEL_ADDR_WIDTH-1 DOWNTO 0)			:= (OTHERS => '1');	
	CONSTANT	MAX_QUADRANT_SIZE			:	STD_LOGIC_VECTOR(QUADRANT_ADDR_WIDTH-1 DOWNTO 0)		:= (OTHERS => '1');	
	CONSTANT	MAX_MAP_SIZE				:	STD_LOGIC_VECTOR(MAP_ADDR_WIDTH-1 DOWNTO 0)				:= (OTHERS => '1');	
	
	--===================================================
	--             MEMORY MAP
	--===================================================
	CONSTANT START_BIT_OFFSET				:	STD_LOGIC_VECTOR(ADDR_AVALON_WIDTH-1 DOWNTO 0) 	:= std_logic_vector(to_unsigned(0,ADDR_AVALON_WIDTH));
	CONSTANT POINTCLOUD_SIZE_OFFSET		:	STD_LOGIC_VECTOR(ADDR_AVALON_WIDTH-1 DOWNTO 0) 	:= std_logic_vector(to_unsigned(1,ADDR_AVALON_WIDTH));
	CONSTANT SIN_THETA_OFFSET				:	STD_LOGIC_VECTOR(ADDR_AVALON_WIDTH-1 DOWNTO 0) 	:= std_logic_vector(to_unsigned(2,ADDR_AVALON_WIDTH));
	CONSTANT COS_THETA_OFFSET				:	STD_LOGIC_VECTOR(ADDR_AVALON_WIDTH-1 DOWNTO 0) 	:= std_logic_vector(to_unsigned(3,ADDR_AVALON_WIDTH));
	CONSTANT DIFF_X_OFFSET					:	STD_LOGIC_VECTOR(ADDR_AVALON_WIDTH-1 DOWNTO 0) 	:= std_logic_vector(to_unsigned(4,ADDR_AVALON_WIDTH));
	CONSTANT DIFF_Y_OFFSET					:	STD_LOGIC_VECTOR(ADDR_AVALON_WIDTH-1 DOWNTO 0) 	:= std_logic_vector(to_unsigned(5,ADDR_AVALON_WIDTH));
	CONSTANT DONE_TICK_OFFSET				:	STD_LOGIC_VECTOR(ADDR_AVALON_WIDTH-1 DOWNTO 0) 	:= std_logic_vector(to_unsigned(6,ADDR_AVALON_WIDTH));
	CONSTANT MAP_SIZE_REG_OFFSET			:	STD_LOGIC_VECTOR(ADDR_AVALON_WIDTH-1 DOWNTO 0) 	:= std_logic_vector(to_unsigned(7,ADDR_AVALON_WIDTH));
	CONSTANT UPDATE_VALID					:	STD_LOGIC_VECTOR(ADDR_AVALON_WIDTH-1 DOWNTO 0) 	:= std_logic_vector(to_unsigned(8,ADDR_AVALON_WIDTH));
	CONSTANT INPUT_DATA_OFFSET				:	STD_LOGIC_VECTOR(ADDR_AVALON_WIDTH-1 DOWNTO 0) 	:= std_logic_vector(to_unsigned(9,ADDR_AVALON_WIDTH));
	CONSTANT INPUT_DATA_OFFSET_UNSIGNED	:	UNSIGNED(ADDR_AVALON_WIDTH-1 DOWNTO 0) 			:= to_unsigned(9,ADDR_AVALON_WIDTH);
	CONSTANT OUTPUT_DATA_OFFSET			:	STD_LOGIC_VECTOR(ADDR_AVALON_WIDTH-1 DOWNTO 0) 	:= std_logic_vector(to_unsigned(16394,ADDR_AVALON_WIDTH));
	CONSTANT OUTPUT_DATA_OFFSET_UNSIGNED:	UNSIGNED(ADDR_AVALON_WIDTH-1 DOWNTO 0) 			:= to_unsigned(16394,ADDR_AVALON_WIDTH);

	CONSTANT	X_LSB								:	INTEGER														:= 0;
	CONSTANT	X_MSB								:	INTEGER														:= 31;
	CONSTANT	Y_LSB								:	INTEGER														:= 32;
	CONSTANT	Y_MSB								:	INTEGER														:= 63;
	CONSTANT	Z_LSB								:	INTEGER														:= 64;
	CONSTANT	Z_MSB								:	INTEGER														:= 95;
	
	
	--===================================================
	--             TYPE DECLARATIONS
	--===================================================
	--type quadrant_memory IS ARRAY(natural range <>) OF STD_LOGIC_VECTOR;
	--type quadrant_memory IS ARRAY(0 to 15) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
	
	
	
END PACKAGE my_package;

	
	
